-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Nov 03 21:15:22 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ST_MACH IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC
    );
END ST_MACH;

ARCHITECTURE BEHAVIOR OF ST_MACH IS
    TYPE type_fstate IS (A,B,C,D);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_z : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x,reg_z)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            reg_z <= '0';
            z <= '0';
        ELSE
            reg_z <= '0';
            z <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '0')) THEN
                        reg_fstate <= B;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    IF ((x = '1')) THEN
                        reg_z <= '1';
                    ELSIF ((x = '0')) THEN
                        reg_z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_z <= '0';
                    END IF;
                WHEN B =>
                    IF ((x = '1')) THEN
                        reg_fstate <= A;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;

                    IF ((x = '0')) THEN
                        reg_z <= '0';
                    ELSIF ((x = '1')) THEN
                        reg_z <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_z <= '0';
                    END IF;
                WHEN C =>
                    IF ((x = '0')) THEN
                        reg_fstate <= D;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    IF ((x = '0')) THEN
                        reg_z <= '1';
                    ELSIF ((x = '1')) THEN
                        reg_z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_z <= '0';
                    END IF;
                WHEN D =>
                    IF ((x = '1')) THEN
                        reg_fstate <= A;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= D;
                    END IF;

                    IF ((x = '0')) THEN
                        reg_z <= '0';
                    ELSIF ((x = '1')) THEN
                        reg_z <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_z <= '0';
                    END IF;
                WHEN OTHERS => 
                    reg_z <= 'X';
                    report "Reach undefined state";
            END CASE;
            z <= reg_z;
        END IF;
    END PROCESS;
END BEHAVIOR;
